library IEEE;
use IEEE.std_logic_1164.all;

entity memory_hierarchy is
  port(
    instruction_cache_data    : in  std_logic_vector(31 downto 0);
    instruction_cache_address : in  std_logic_vector(31 downto 0);
    data_cache_data           : in  std_logic_vector(31 downto 0);
    data_cache_address        : in  std_logic_vector(31 downto 0);
    RW                        : in  std_logic;
    clk                       : in  std_logic;
    ready                     : out std_logic
    );
end entity;

architecture arch of memory_hierarchy is

component control_unit is
  port(
    RW                      : in  std_logic;
    enable                  : in  std_logic;
    buffer_ready            : in  std_logic;
    data_cache_ready        : in  std_logic;
    instruction_cache_ready : in  std_logic;
    data_cache_hit          : in  boolean;
    instruction_cache_hit   : in  boolean;
    clk                     : in  std_logic;  -- clock de periodo 5 ns
    SEL                     : out std_logic_vector(1 downto 0);
    ready                   : out std_logic
    );
end component;

component instruction_cache is
  port (
    data    : out std_logic_vector(31 downto 0);
    address : in  std_logic_vector(31 downto 0);
    enable  : in  std_logic;
    ready   : out std_logic;
    hit: out boolean;
    clk     : in  std_logic
    );
end component;

component data_cache is
  port (
    data_in  : in  std_logic_vector(31 downto 0);
    data_out : out std_logic_vector(31 downto 0);
    ADDR32   : in  std_logic_vector(31 downto 0);
    RW       : in  std_logic;           -- 0 para Read, 1 para Write
    ENABLE   : in  std_logic;
    READY    : out std_logic;
    hit      : out boolean;
    clk      : in  std_logic
    );
end component;

component main_memory is
  generic (
    filename   : in string;
    read_time  : in time := 40 ns;
    write_time : in time := 40 ns
    );
  port (
    data    : inout std_logic_vector(31 downto 0);
    address : in    std_logic_vector(31 downto 0);
    rw      : in    std_logic;
    enable  : in    std_logic;
    ready   : out   std_logic
    );
end component;

begin
end arch;
